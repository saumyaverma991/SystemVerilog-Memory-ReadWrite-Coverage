// Code your testbench here
// or browse Examples
/*typedef class monitor;
typedef class generator;
typedef class coverage;
typedef class agent;
typedef class common;
typedef class bfm;
typedef class env;
typedef class tx;
*/
`include "common_c.sv"
`include "interface_c.sv"
`include "transaction_c.sv"
`include "generator_c.sv"
`include "bfm_c.sv"
`include "coverage_c.sv"
`include "monitor_c.sv"
`include "agent_c.sv"
`include "environment_c.sv"
`include "memory.sv"
`include "top_c.sv"


